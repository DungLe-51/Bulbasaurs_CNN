module conv_layer #(

)(

);
endmodule